** Profile: "SCHEMATIC1-Worst_Case"  [ D:\Orcad Work\cdssetup\workspace\projects\draft_proiect_paul\draft_proiect_paul-pspicefiles\schematic1\worst_case.sim ] 

** Creating circuit file "Worst_Case.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Orcad Work/cdssetup/workspace/projects/draft_proiect2/diodaled.lib" 
* From [PSPICE NETLIST] section of D:\Orcad Work\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 10u 
.WCASE TRAN V([OUT]) YMAX VARY BOTH  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
