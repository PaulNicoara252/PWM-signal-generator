** Profile: "SCHEMATIC1-dioda"  [ D:\Orcad Work\cdssetup\workspace\projects\draft_proiect_paul\Draft_proiect_PAUL-PSpiceFiles\SCHEMATIC1\dioda.sim ] 

** Creating circuit file "dioda.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Orcad Work/cdssetup/workspace/projects/draft_proiect2/diodaled.lib" 
* From [PSPICE NETLIST] section of D:\Orcad Work\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V3 0 5 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
