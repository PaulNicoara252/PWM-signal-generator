** Profile: "SCHEMATIC1-Parametric_Sweep"  [ D:\Orcad Work\cdssetup\workspace\projects\draft_proiect_paul\draft_proiect_paul-pspicefiles\schematic1\parametric_sweep.sim ] 

** Creating circuit file "Parametric_Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Orcad Work/cdssetup/workspace/projects/draft_proiect2/diodaled.lib" 
* From [PSPICE NETLIST] section of D:\Orcad Work\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.25m 0 
.STEP LIN PARAM cursor1 0 1 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
