** Profile: "SCHEMATIC1-Analiza_Monte_Carlo"  [ D:\Orcad Work\cdssetup\workspace\projects\draft_proiect_paul\draft_proiect_paul-pspicefiles\schematic1\analiza_monte_carlo.sim ] 

** Creating circuit file "Analiza_Monte_Carlo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Orcad Work/cdssetup/workspace/projects/draft_proiect2/diodaled.lib" 
* From [PSPICE NETLIST] section of D:\Orcad Work\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 
.MC 100 TRAN V([OUT]) YMAX OUTPUT ALL 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
